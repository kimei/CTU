kimei@COMPETReadout003.23511:1320922768