LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY system IS
PORT (
	fpga_0_RS232_sin_pin : IN STD_LOGIC;
	fpga_0_RS232_sout_pin : OUT STD_LOGIC;
	fpga_0_LEDs_8Bit_GPIO_d_out_pin : OUT STD_LOGIC_VECTOR(0 TO 7);
	fpga_0_DIP_Switches_8Bit_GPIO_in_pin : IN STD_LOGIC_VECTOR(0 TO 7);
	fpga_0_Push_Buttons_3Bit_GPIO_in_pin : IN STD_LOGIC_VECTOR(0 TO 2);
	fpga_0_FLASH_8Mx16_Mem_DQ_pin : INOUT STD_LOGIC_VECTOR(0 TO 15);
	fpga_0_FLASH_8Mx16_Mem_A_pin : OUT STD_LOGIC_VECTOR(7 TO 31);
	fpga_0_FLASH_8Mx16_Mem_WEN_pin : OUT STD_LOGIC;
	fpga_0_FLASH_8Mx16_Mem_OEN_pin : OUT STD_LOGIC_VECTOR(0 TO 0);
	fpga_0_FLASH_8Mx16_Mem_CEN_pin : OUT STD_LOGIC_VECTOR(0 TO 0);
	fpga_0_FLASH_8Mx16_rpn_dummy_pin : OUT STD_LOGIC;
	fpga_0_FLASH_8Mx16_byte_dummy_pin : OUT STD_LOGIC;
	fpga_0_FLASH_8Mx16_adv_dummy_pin : OUT STD_LOGIC;
	fpga_0_FLASH_8Mx16_clk_dummy_pin : OUT STD_LOGIC;
	fpga_0_FLASH_8Mx16_wait_dummy_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_ODT_pin : OUT STD_LOGIC_VECTOR(0 TO 0);
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_A_pin : OUT STD_LOGIC_VECTOR(12 DOWNTO 0);
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_BA_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_CAS_N_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_CKE_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_CS_N_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_RAS_N_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_WE_N_pin : OUT STD_LOGIC;
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_DM_pin : OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_DQS : INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_DQS_N : INOUT STD_LOGIC_VECTOR(3 DOWNTO 0);
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_DQ : INOUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_CK_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_DDR2_SDRAM_16Mx32_DDR2_CK_N_pin : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
	fpga_0_Hard_Ethernet_MAC_TemacPhy_RST_n_pin : OUT STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_GMII_TXD_0_pin : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
	fpga_0_Hard_Ethernet_MAC_GMII_TX_EN_0_pin : OUT STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_GMII_TX_CLK_0_pin : OUT STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_GMII_TX_ER_0_pin : OUT STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_GMII_RX_ER_0_pin : IN STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_GMII_RX_CLK_0_pin : IN STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_GMII_RX_DV_0_pin : IN STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_GMII_RXD_0_pin : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
	fpga_0_Hard_Ethernet_MAC_MII_TX_CLK_0_pin : IN STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_MDC_0_pin : OUT STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_MDIO_0_pin : INOUT STD_LOGIC;
	fpga_0_Hard_Ethernet_MAC_PHY_MII_INT_pin : OUT STD_LOGIC;
	sys_clk_pin : IN STD_LOGIC;
	sys_rst_pin : IN STD_LOGIC
	);
END system;

ARCHITECTURE STRUCTURE OF system IS

BEGIN
END ARCHITECTURE STRUCTURE;
